Inverter: Basic Example

* Technology Dependent design rules/parameters
.include /CMC/setups/ensc450/HSPICE/cmosp18/rules.inc
* Wm#, Awd# parameters etc. all specified in the rules.inc file above

* Transistor models 
.protect
.LIB `/CMC/setups/ensc450/HSPICE/cmosp18/log018.l' SS  $ typical process corner.
.unprotect

* Supply Sources
.param pwr=1.05 
.temp 125
Vvdd  vdd  0 dc pwr
Vvdds vdds 0 dc pwr
Vgnd  gnd  0 dc 0
Vgnds gnds 0 dc 0

* Logic 
.param Wn=Wm#
Xpmos vdd a z vdds pt_st w=2*Wn
Xnmos gnd a z gnds nt_st w=Wn

Cload z 0 20f

* Input Stimuli (Step response)
VA  a  0 PWL(0n 0 9ns 0 10ns pwr)


* Simulation Parameters ************************
.tran 0.01ps 40ns START=0
* Sweeps transistor width 
* .tran 0.01ps 40ns START=0 sweep Wn START=Wn STOP=4*Wn STEP=Wn 

.graph V(a)
.graph V(z)
.option post

* Measure propogation delay from rising edge of input A to falling edge of output Z
.meas tran tpd_in01      trig v(a) val='pwr*0.5' cross=1
+                        targ v(z) val='pwr*0.5' cross=1 

* Measure output delay from falling edge of output Z
.meas tran ttr           trig v(z) val='pwr*0.8' fall=1
+                        targ v(z) val='pwr*0.2' fall=1

* Measures Power (cell leakage and dynamic)
.meas tran leak_pow_in1  avg power FROM=12ns TO=14ns
.meas tran leak_pow_in0  avg power FROM= 6ns TO= 8ns
.meas tran dyn_pow       avg power FROM= 9ns TO=10ns

************************************************

.end
  
